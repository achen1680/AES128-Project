module add_roundkey(

);